library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;
entity rom_memory is
    Port ( addr : in STD_LOGIC_VECTOR (10 downto 0);
           dout_curr : out STD_LOGIC_VECTOR (31 downto 0);
           dout_prev : out STD_LOGIC_VECTOR (31 downto 0));
end rom_memory;

architecture Behavioral of rom_memory is

type matrix is array(0 to 1700) of integer;

signal content: matrix := (
    2734,
    2100,
    4688,
    2344,
    3027,
    3906,
    2148,
    2393,
    4346,
    2100,
    2295,
    2686,
    4541,
    2295,
    2393,
    4150,
    2344,
    2100,
    2051,
    2051,
    3857,
    2295,
    2246,
    2148,
    4395,
    2344,
    4541,
    3564,
    2051,
    4639,
    3760,
    4688,
    2197,
    2148,
    2295,
    4395,
    2197,
    2197,
    2295,
    4443,
    2148,
    2002,
    3613,
    2148,
    2100,
    2002,
    2100,
    2441,
    2246,
    2051,
    3271,
    2637,
    2148,
    3661,
    2637,
    2100,
    2148,
    4590,
    4199,
    3515,
    2148,
    3125,
    2051,
    2637,
    4785,
    2051,
    3271,
    4492,
    2051,
    3174,
    2490,
    3076,
    3076,
    3760,
    3076,
    3515,
    2051,
    2148,
    2441,
    4248,
    3809,
    2539,
    2246,
    2002,
    3661,
    4346,
    3271,
    2002,
    2002,
    3661,
    2930,
    2002,
    2246,
    2246,
    2002,
    2197,
    2148,
    2051,
    3954,
    2100,
    2344,
    3661,
    4346,
    2441,
    2197,
    3711,
    4639,
    2051,
    1953,
    2100,
    2100,
    2002,
    2637,
    3564,
    3320,
    3661,
    2148,
    2051,
    2783,
    2002,
    4590,
    2148,
    4150,
    4004,
    2148,
    2002,
    3906,
    2051,
    2002,
    2051,
    2344,
    2002,
    4395,
    2051,
    3320,
    4736,
    3418,
    3125,
    3711,
    2051,
    4150,
    2344,
    2588,
    2051,
    2148,
    2881,
    4150,
    2148,
    2051,
    2051,
    2246,
    4199,
    2490,
    2051,
    2246,
    2148,
    2441,
    2295,
    2051,
    2246,
    2441,
    2441,
    4736,
    2295,
    2100,
    2539,
    2197,
    2197,
    2393,
    2295,
    3222,
    4102,
    3320,
    3613,
    2197,
    2100,
    2246,
    2441,
    3760,
    2734,
    2197,
    2246,
    2441,
    2295,
    2588,
    2148,
    2197,
    3125,
    2148,
    3467,
    2539,
    2197,
    4492,
    2637,
    2979,
    2979,
    3857,
    2246,
    3222,
    2148,
    4541,
    2393,
    4639,
    2344,
    3613,
    2441,
    4443,
    2637,
    3271,
    3369,
    2148,
    2734,
    3711,
    2148,
    3906,
    2832,
    2246,
    2295,
    3467,
    3027,
    2588,
    2637,
    4492,
    2246,
    3320,
    2295,
    2246,
    3906,
    4492,
    4443,
    2295,
    3711,
    2588,
    3613,
    2295,
    2490,
    3467,
    2637,
    2490,
    2246,
    4639,
    2246,
    2246,
    3564,
    2246,
    2539,
    2393,
    2588,
    3369,
    2246,
    2246,
    2295,
    3027,
    3467,
    2344,
    2246,
    4395,
    2344,
    2637,
    2246,
    2295,
    2246,
    3271,
    2441,
    3369,
    2246,
    2246,
    2637,
    2246,
    4102,
    2344,
    2295,
    2246,
    2588,
    3467,
    4443,
    3125,
    4248,
    2295,
    2539,
    4102,
    3613,
    3661,
    2295,
    2246,
    4248,
    2832,
    3369,
    2344,
    2344,
    2588,
    2295,
    3125,
    2490,
    2246,
    2295,
    4150,
    3467,
    2734,
    2734,
    2686,
    2441,
    2539,
    4346,
    2441,
    2539,
    2490,
    4395,
    3906,
    2441,
    3954,
    4395,
    3467,
    2588,
    2393,
    3711,
    2539,
    3515,
    2539,
    2295,
    2295,
    4346,
    2344,
    2393,
    2539,
    2539,
    2441,
    4541,
    3320,
    2734,
    2246,
    4541,
    2832,
    2588,
    2295,
    3271,
    3222,
    2246,
    3711,
    2246,
    3418,
    4541,
    4150,
    2441,
    2539,
    2930,
    4004,
    2637,
    2539,
    2637,
    4639,
    2686,
    2344,
    2686,
    2344,
    2686,
    2539,
    3564,
    4248,
    4541,
    3906,
    3711,
    2588,
    2295,
    3564,
    2686,
    4395,
    3418,
    2295,
    2246,
    2490,
    2344,
    2441,
    2393,
    2686,
    3125,
    2637,
    2686,
    3369,
    2734,
    3809,
    2832,
    2441,
    2295,
    2295,
    2393,
    2539,
    2588,
    2686,
    2930,
    2393,
    2441,
    2783,
    2686,
    2295,
    2344,
    2686,
    3369,
    3174,
    3661,
    3809,
    2295,
    2344,
    2832,
    2734,
    2441,
    3467,
    2686,
    2393,
    2734,
    2490,
    2490,
    3271,
    4346,
    2295,
    2734,
    2295,
    2295,
    4492,
    3418,
    2588,
    2539,
    3125,
    2783,
    4395,
    2539,
    2393,
    2344,
    3661,
    2344,
    2490,
    2344,
    2588,
    2734,
    2344,
    2588,
    2295,
    2441,
    4199,
    2930,
    2295,
    2246,
    4639,
    4395,
    2295,
    2246,
    3954,
    3027,
    3320,
    2441,
    3857,
    4590,
    4346,
    3809,
    3954,
    2734,
    2295,
    3760,
    2246,
    3174,
    2441,
    4395,
    3076,
    2686,
    2344,
    3076,
    3467,
    4492,
    2930,
    2539,
    2393,
    2490,
    2393,
    2832,
    2295,
    3320,
    2295,
    2539,
    2295,
    3515,
    2393,
    3613,
    2246,
    2246,
    2393,
    2539,
    4150,
    3174,
    4346,
    2539,
    2295,
    2539,
    2637,
    2539,
    4297,
    2881,
    2734,
    3027,
    2441,
    2930,
    4248,
    3320,
    2295,
    2295,
    3661,
    2637,
    4199,
    2246,
    2295,
    4346,
    3760,
    2295,
    4150,
    2246,
    2686,
    4297,
    2393,
    3076,
    2441,
    2734,
    2539,
    2344,
    2734,
    2734,
    2490,
    2930,
    2832,
    2490,
    3711,
    3515,
    2197,
    2295,
    2637,
    4688,
    4541,
    2686,
    2344,
    2783,
    3467,
    2344,
    4297,
    3954,
    2344,
    2441,
    4053,
    2979,
    2979,
    2979,
    2979,
    2979,
    2979,
    2979,
    2979,
    2979,
    3027,
    2979,
    2979,
    2979,
    3027,
    3027,
    2979,
    3027,
    3027,
    3027,
    3027,
    3027,
    3027,
    3027,
    3027,
    3076,
    3076,
    3076,
    3027,
    3027,
    3076,
    3076,
    3027,
    3076,
    3076,
    3076,
    3027,
    3027,
    3027,
    3076,
    3076,
    3076,
    3076,
    3076,
    3076,
    3076,
    3076,
    3076,
    2832,
    3125,
    2588,
    2588,
    2734,
    2734,
    2783,
    3222,
    3174,
    4541,
    2832,
    3174,
    2734,
    2637,
    4297,
    3027,
    2881,
    2979,
    2930,
    3515,
    4932,
    4541,
    3125,
    2783,
    2686,
    3564,
    2588,
    2637,
    2588,
    3760,
    2637,
    4150,
    2637,
    2686,
    3711,
    2734,
    2686,
    2686,
    2832,
    3076,
    3125,
    2637,
    2832,
    3174,
    4297,
    3711,
    4346,
    3271,
    4297,
    2734,
    3125,
    4639,
    2783,
    2734,
    3027,
    4834,
    4785,
    2734,
    3760,
    4102,
    3222,
    3125,
    2881,
    2881,
    3174,
    2979,
    3661,
    2881,
    3125,
    2881,
    4102,
    3857,
    4395,
    3467,
    2783,
    3222,
    2881,
    3174,
    2930,
    3369,
    4492,
    2930,
    2930,
    2930,
    3369,
    3125,
    3271,
    3418,
    3320,
    3369,
    3125,
    4199,
    2979,
    3320,
    3369,
    3271,
    3076,
    3418,
    4980,
    3515,
    3222,
    4883,
    3174,
    3467,
    3564,
    3613,
    3613,
    3222,
    3564,
    3222,
    3271,
    3954,
    3174,
    3564,
    3711,
    3613,
    4004,
    3271,
    4248,
    3271,
    3076,
    4443,
    3369,
    3613,
    4639,
    2832,
    3418,
    2783,
    3027,
    3320,
    3271,
    3613,
    2832,
    2979,
    3027,
    3174,
    3954,
    3369,
    3125,
    3174,
    3369,
    3125,
    3076,
    4102,
    2832,
    2930,
    2783,
    3174,
    2832,
    3174,
    3222,
    3369,
    2734,
    3271,
    3467,
    3613,
    2783,
    3369,
    3027,
    2979,
    2832,
    3222,
    3369,
    2783,
    2783,
    3320,
    2832,
    2930,
    2783,
    3271,
    2832,
    2783,
    3760,
    3515,
    3369,
    3222,
    3271,
    3027,
    3906,
    3076,
    3271,
    2979,
    4004,
    3125,
    3174,
    3857,
    3222,
    4443,
    3076,
    3174,
    2881,
    3271,
    3125,
    3125,
    3076,
    3125,
    3125,
    2832,
    3418,
    2930,
    2979,
    3271,
    3125,
    2881,
    2832,
    4053,
    2930,
    3271,
    2930,
    2832,
    3174,
    4443,
    4492,
    2832,
    2881,
    3320,
    4053,
    3222,
    3369,
    2832,
    4639,
    2832,
    3076,
    2881,
    2979,
    3857,
    2881,
    4443,
    3418,
    3320,
    4590,
    3027,
    3174,
    4590,
    2881,
    2881,
    3076,
    2881,
    4053,
    3369,
    3125,
    3369,
    3320,
    3076,
    4541,
    2881,
    3320,
    3222,
    2930,
    2832,
    3174,
    3515,
    2832,
    4639,
    2832,
    2930,
    4346,
    2930,
    2930,
    3125,
    3369,
    2832,
    4639,
    2930,
    3027,
    2881,
    3661,
    3076,
    3027,
    3954,
    3613,
    3076,
    3369,
    4346,
    3760,
    3125,
    3076,
    4053,
    2930,
    3222,
    3711,
    3222,
    3369,
    4346,
    3222,
    2930,
    3906,
    3467,
    3320,
    3418,
    4150,
    3809,
    3125,
    4150,
    4297,
    3027,
    3564,
    3125,
    2930,
    3271,
    3027,
    3271,
    3174,
    3564,
    3564,
    4102,
    3320,
    3174,
    3320,
    3467,
    3271,
    3174,
    3711,
    3125,
    3467,
    3222,
    4590,
    4248,
    3320,
    3369,
    3222,
    4297,
    3222,
    3125,
    3174,
    3174,
    4199,
    3661,
    4102,
    3661,
    3222,
    3125,
    3613,
    3467,
    3271,
    3613,
    3711,
    3174,
    3515,
    4297,
    4395,
    3174,
    3661,
    3418,
    3222,
    3418,
    4492,
    4102,
    3515,
    3613,
    3857,
    3320,
    3467,
    3467,
    3809,
    4443,
    3125,
    3661,
    3271,
    3125,
    3564,
    3515,
    4541,
    4004,
    3125,
    3125,
    4590,
    3125,
    3174,
    3613,
    3564,
    3467,
    3613,
    3125,
    3369,
    4443,
    3320,
    3125,
    3125,
    3418,
    4541,
    3320,
    3320,
    3222,
    4053,
    3418,
    3564,
    3564,
    3369,
    3125,
    3125,
    3661,
    3320,
    4346,
    3174,
    3613,
    3661,
    4297,
    3076,
    4590,
    3174,
    3271,
    3271,
    3418,
    3174,
    3613,
    4102,
    3369,
    3418,
    3271,
    3320,
    3076,
    3613,
    3222,
    4395,
    3076,
    4395,
    3076,
    4199,
    3222,
    3711,
    3661,
    3369,
    3954,
    3906,
    3564,
    3613,
    3418,
    3613,
    3369,
    3125,
    3174,
    3125,
    3125,
    3125,
    4346,
    4004,
    4395,
    3418,
    3809,
    3467,
    3661,
    3125,
    3125,
    3174,
    3174,
    3711,
    3125,
    3661,
    3125,
    3564,
    3320,
    3125,
    3906,
    3613,
    3125,
    3320,
    3125,
    3613,
    3222,
    3613,
    3222,
    4541,
    3271,
    3515,
    3857,
    3564,
    3613,
    3320,
    3857,
    3467,
    4395,
    3320,
    3174,
    3320,
    3564,
    3564,
    3125,
    3125,
    3125,
    3369,
    3125,
    3418,
    4346,
    3125,
    3515,
    3613,
    3174,
    3125,
    4346,
    3271,
    3613,
    3320,
    3125,
    3418,
    3809,
    3613,
    3369,
    3613,
    3125,
    3125,
    3222,
    4248,
    3125,
    3711,
    3174,
    4443,
    3711,
    3174,
    3564,
    3711,
    3222,
    4150,
    3271,
    3320,
    3369,
    3613,
    3613,
    3760,
    4492,
    3174,
    3954,
    3174,
    3711,
    3320,
    3222,
    3515,
    3711,
    4297,
    3564,
    3271,
    3174,
    4053,
    3613,
    3271,
    3174,
    3857,
    3418,
    3222,
    3760,
    3271,
    3515,
    3809,
    3320,
    3174,
    3564,
    3954,
    3954,
    3418,
    3369,
    3954,
    3222,
    3418,
    3954,
    3467,
    3467,
    4297,
    3760,
    3613,
    3467,
    4053,
    3369,
    3906,
    4541,
    3271,
    3271,
    3564,
    3467,
    3369,
    3418,
    3467,
    3661,
    4102,
    3760,
    3661,
    3661,
    3661,
    3613,
    3174,
    3222,
    4199,
    3711,
    3467,
    3320,
    3222,
    3222,
    3467,
    3271,
    3369,
    3222,
    3564,
    3760,
    3711,
    4150,
    3222,
    3613,
    3467,
    3613,
    3320,
    3467,
    4492,
    3222,
    3564,
    3613,
    3564,
    3467,
    4541,
    3320,
    3369,
    3320,
    3369,
    3467,
    3369,
    3467,
    3857,
    3271,
    3467,
    3515,
    3760,
    3174,
    3418,
    3613,
    3954,
    3613,
    3857,
    3174,
    3271,
    3125,
    3271,
    3418,
    3467,
    3174,
    3174,
    3174,
    3222,
    3174,
    4492,
    3222,
    4102,
    3418,
    3271,
    3418,
    3711,
    3222,
    3320,
    3661,
    4102,
    3222,
    3222,
    3613,
    3222,
    3661,
    4395,
    3711,
    3271,
    3564,
    3174,
    3711,
    3174,
    3320,
    4443,
    3711,
    3369,
    3857,
    3222,
    4297,
    3467,
    3418,
    3271,
    4102,
    3418,
    4199,
    4004,
    3418,
    3222,
    3515,
    3711,
    3418,
    3271,
    3369,
    3515,
    3760,
    3222,
    3174,
    4199,
    3515,
    4053,
    3711,
    3271,
    4297,
    4053,
    3613,
    3174,
    3613,
    3271,
    3418,
    4297,
    3418,
    3661,
    3857,
    3467,
    4053,
    3613,
    3174,
    3125,
    3661,
    3809,
    3515,
    4541,
    3418,
    3271,
    3125,
    3418,
    3320,
    3320,
    3515,
    4004,
    4102,
    3564,
    3711,
    3174,
    3564,
    4102,
    3711,
    3320,
    3515,
    3369,
    3222,
    3564,
    3711,
    3320,
    3857,
    3711,
    3760,
    3320,
    3174,
    3564,
    3125,
    3174,
    3661,
    3174,
    3418,
    3369,
    3711,
    3418,
    3222,
    3418,
    3857,
    3515,
    3906,
    3857,
    3222,
    3320,
    4004,
    3661,
    3369,
    3222,
    3125,
    4443,
    3174,
    3125,
    3125,
    3760,
    3125,
    3174,
    3661,
    3809,
    3174,
    3613,
    3320,
    3613,
    3369,
    3515,
    3613,
    3174,
    4004,
    3125,
    3320,
    3125,
    3174,
    3418,
    3613,
    4443,
    3125,
    3613,
    3369,
    3125,
    3467,
    3613,
    3320,
    3418,
    3222,
    3515,
    3174,
    3369,
    3564,
    3222,
    4443,
    3271,
    3906,
    3467,
    3418,
    3174,
    4443,
    3076,
    3369,
    4297,
    3760,
    3613,
    3369,
    3125,
    3661,
    3564,
    3857,
    3857,
    3222,
    3320,
    3906,
    3661,
    3369,
    3369,
    3711,
    3076,
    3076,
    3125,
    3515,
    3320,
    3564,
    3564,
    3320,
    3174,
    3613,
    3076,
    3222,
    3174,
    3467,
    3613,
    3564,
    3760,
    4395,
    3369,
    3515,
    3613,
    3222,
    3613,
    3174,
    3125,
    3125,
    3418,
    3125,
    3418,
    3222,
    3661,
    3564,
    3222,
    3125,
    3711,
    3564,
    3711,
    3320,
    3564,
    3857,
    3271,
    3320,
    3125,
    3760,
    3222,
    3515,
    3320,
    3369,
    3271,
    3760,
    4639,
    3320,
    3222,
    3661,
    3760,
    3760,
    3661,
    3515,
    3564,
    4199,
    3222,
    3271,
    4590,
    3174,
    3174,
    3564,
    3809,
    3467,
    3515,
    3271,
    3954,
    3174,
    4395,
    3222,
    3369,
    3174,
    3564,
    3271,
    3271,
    3613,
    4004,
    3809,
    3174,
    3369,
    3369,
    3271,
    3222,
    4736,
    3711,
    3760,
    4688,
    3320,
    3809,
    4297,
    3271,
    3222,
    3320,
    4639,
    3320,
    3174,
    3418,
    3222,
    3271,
    4785,
    3222,
    3711,
    4834,
    3467,
    3760,
    3467,
    4932,
    3174,
    3613,
    3369,
    3271,
    3515,
    3222,
    3515,
    3760,
    3661,
    3661,
    3711,
    3515,
    3369,
    3564,
    3418,
    3564,
    3271,
    3809,
    3467,
    3271,
    3857,
    3760,
    4395,
    3711,
    3418,
    3271,
    4590,
    3320,
    3222,
    3320,
    3515,
    3613,
    3418,
    3857,
    3222,
    3661,
    3564,
    3515,
    3906,
    3760,
    3906,
    3320,
    4395,
    3809,
    4932,
    3320,
    3564,
    3320,
    4492,
    3467,
    3369,
    4199,
    3613,
    3564,
    3418,
    3369,
    4492,
    3418,
    3369,
    4590,
    3418,
    3906,
    3613,
    3711,
    3467,
    3515,
    3467,
    4053,
    4834,
    3564,
    3467,
    3613,
    3857,
    3954,
    3613,
    3809,
    4541,
    3418,
    3711,
    3809,
    4688,
    3418,
    3418,
    3906,
    3613,
    4395,
    3613,
    3613,
    4932,
    3661,
    3467,
    3369,
    3613,
    3418,
    4541,
    3320,
    3661,
    3418,
    3760,
    3857,
    3320,
    3320,
    3661,
    3418,
    3661,
    3906,
    3564,
    4883,
    3711,
    3515,
    3271,
    3369,
    3613,
    3320,
    4443,
    3271,
    3320,
    3857,
    4395,
    4639,
    3857,
    3857,
    3418,
    3809,
    3369,
    3760,
    3809,
    3320,
    3369,
    3906,
    3564,
    3906,
    4199,
    3661,
    3467,
    4639,
    3369,
    3661,
    4590,
    3564,
    4004,
    3418,
    3320,
    3369,
    3515,
    3906,
    3515,
    4590,
    3711,
    4395,
    3418,
    3613,
    3661,
    3320,
    3613,
    3857,
    3613,
    3418,
    3564,
    3467,
    4492,
    3467,
    3320,
    4004,
    3760,
    3613,
    3857,
    4199,
    3467,
    4541,
    4297,
    3954,
    4541,
    3320,
    3271,
    3320
);
begin

    dout_curr <= std_logic_vector(to_signed(content(to_integer(unsigned(addr))), 32));
    dout_prev <= std_logic_vector(to_signed(content(to_integer(unsigned(addr - 1))), 32));

end Behavioral;